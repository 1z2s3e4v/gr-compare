version https://git-lfs.github.com/spec/v1
oid sha256:42b26779263fca144c55703e28353c5038a768d4478caf442f45d3fde75fba01
size 299111
