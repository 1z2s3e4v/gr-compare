version https://git-lfs.github.com/spec/v1
oid sha256:ec9d9376d979a90cb5b12b75a27d7fd98770bb48fafaeccfa448fc7f47b00ca6
size 284656
