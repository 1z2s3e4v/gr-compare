version https://git-lfs.github.com/spec/v1
oid sha256:558e1e7387505c405715ca0b14a4b063f525bea31fd0ab496150bae01edc687e
size 196996
