version https://git-lfs.github.com/spec/v1
oid sha256:80a6219a9f9be0b8f6f39cf3dcc49e958280736a111416047495b15bf2d70e57
size 721588
