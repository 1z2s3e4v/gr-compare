version https://git-lfs.github.com/spec/v1
oid sha256:995163295c1365367a3ab07bfba990edda81e8af368074a56dd5ef0ea0cc4355
size 269031
