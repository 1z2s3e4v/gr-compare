version https://git-lfs.github.com/spec/v1
oid sha256:8fefa41b77cd0f15e713e1aa8b541cf7ecf958323210af527fd3715e267e6d58
size 180603
