version https://git-lfs.github.com/spec/v1
oid sha256:88e17b56280c37d766f47ed0a51a8fd984cdebaa1511f03cfe33819834309fb3
size 480622
