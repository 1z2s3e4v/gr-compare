version https://git-lfs.github.com/spec/v1
oid sha256:d50b94524d57e21899a6ec0de049f58d53db56c1f42793f663957cd1db86113f
size 321928
