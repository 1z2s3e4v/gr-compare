version https://git-lfs.github.com/spec/v1
oid sha256:55afc5b234891a3a402f2c8a76d6dac05bfde62457b5dbebf8ccd7568c0d2ab5
size 183336
