version https://git-lfs.github.com/spec/v1
oid sha256:e28d313dc139fe65165b9e756f7b12ae053434a5e62d3a7e24d7507ac6006c44
size 250123
