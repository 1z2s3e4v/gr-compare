version https://git-lfs.github.com/spec/v1
oid sha256:9031a8fccc233b01460de0cf14e9641e40865c3a8bb2d0f390cfe972b24b003e
size 638256
