version https://git-lfs.github.com/spec/v1
oid sha256:bb8fefb913a6cfa28e3dbf606bef791dc01c118b2d284fd97d32cf5ec4f13ec3
size 321699
