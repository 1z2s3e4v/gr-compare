version https://git-lfs.github.com/spec/v1
oid sha256:64f689bab004147c46c6a5cc1fed08303b6e01fbe31755d4f967323aa93354ee
size 270973
