version https://git-lfs.github.com/spec/v1
oid sha256:8c5b90b5e735e751332027c29f3e167a766bf687e1c85b45e46e1f7b71747bdf
size 194286
