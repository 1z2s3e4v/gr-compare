version https://git-lfs.github.com/spec/v1
oid sha256:9e5614e88cea5d50226d76add93af33c459007a4f72122228916beffe2e15af6
size 185617
