version https://git-lfs.github.com/spec/v1
oid sha256:70bf84913ffecba1ffd20242a32d5bb95443c34ba054d3f8f4188973af115f24
size 723311
