version https://git-lfs.github.com/spec/v1
oid sha256:7660a3586715137f5acc10fdbe83e12f3e2e52d8d6d4f7e7ef88b899bec5f03a
size 283636
