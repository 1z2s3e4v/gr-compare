version https://git-lfs.github.com/spec/v1
oid sha256:99cb86b809bcdc332963d965da7a26a1be5907f1a532ce3f06d6370397f487de
size 183313
