version https://git-lfs.github.com/spec/v1
oid sha256:f710bc3c947791e067b4282021a805136477aa5135987ef1280fa414669b6a31
size 287898
