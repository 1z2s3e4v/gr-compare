version https://git-lfs.github.com/spec/v1
oid sha256:674b120641451d26f1051cc62fc1b96cde42addb00841cd3c9b142a064d981f1
size 194286
