version https://git-lfs.github.com/spec/v1
oid sha256:947a047a2acce6eeef50709461e4e5d4455d3f3b9e84a52b3fff034246ea367d
size 723308
