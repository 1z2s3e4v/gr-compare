version https://git-lfs.github.com/spec/v1
oid sha256:087207ea1e3b1a69c801faf4acedd5c1dee1f23a18245c5974ee28690ba5531e
size 795524
